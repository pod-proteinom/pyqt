LOGIC_SW.CIR - BASIC LOGIC GATES USING SWITCHES
*
VCC	10	0	5V
*
* INPUT A AND B, COUNT IN BINARY 0 - 3
VA	1	0	PULSE(5V 0V 0NS 10NS 10NS 90NS 200NS)
VB	2	0	PULSE(5V 0V 0NS 10NS 10NS 190NS 400NS)
*
XNAND1	1 2 3 10	NAND
*
*
* LOGIC GATE SUBCIRCUITS ******************************************
*
.SUBCKT NAND 1 2 3 4
* TERMINALS A B OUT VCC
RL	3	4	500
S1	3 5	1 0 	SW
S2	5 0	2 0 	SW
.ENDS
*
.SUBCKT AND 1 2 3 4
* TERMINALS A B OUT VCC
S1	4 5	1 0 	SW
S2	5 3	2 0 	SW
RL	3	0	500
.ENDS
*
.SUBCKT NOR 1 2 3 4
* TERMINALS A B OUT VCC
RL	3	4	500
S1	3 0	1 0 	SW
S2	3 0	2 0 	SW
.ENDS
*
.SUBCKT NOT 1 3 4
* TERMINALS A OUT VCC
RL	3	4	500
S1	3 0	1 0 	SW
.ENDS
*
*
.MODEL	SW	VSWITCH(VON=2.6 VOFF=2.4 RON=10 ROFF=1MEG)
*
* ANALYSIS **************************************************
.TRAN 	5NS  	400NS
*
* VIEW RESULTS
.PRINT	TRAN 	V(1) V(2) V(3)
.PROBE
.END