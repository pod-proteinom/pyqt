* Adder - 4 bit all-nand-gate binary adder
.SUBCKT NAND 1 2 3 4
* TERMINALS A B OUT VCC
RL	3	4	500
S1	3 5	1 0 	SW
S2	5 0	2 0 	SW
.ENDS

.SUBCKT onearg one
.ENDS

.SUBCKT twoarg one two
.ENDS

.SUBCKT NOT 1 3 4
* TERMINALS A OUT VCC
RL	3	4	500
S1	3 0	1 0 	SW
.ENDS

.subckt ONEBIT 1 2 3 4 5  6
X1 1 2 7 6 NAND
X2 1 7 8 6 NAND
X3 2 7 9 6 NAND
X4 8 9 10 6 NAND
X5 3 10 11 6 NAND
X6 3 11 12 6 NAND
X7 10 11 13 6 NAND
X8 12 13 4 6 NAND
X9 11 7 5 6 NAND
.ends
*
.SUBCKT FOURBIT 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
X1 1 2 13 9 16 15 ONEBIT
X2 3 4 16 10 17 15 ONEBIT
X3 5 6 17 11 18 15 ONEBIT
X4 7 8 18 12 14 15 ONEBIT
.ENDS